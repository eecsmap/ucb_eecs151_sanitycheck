module z1top(
    input BUTTON,
    output LED
);

    assign LED = BUTTON;

endmodule
